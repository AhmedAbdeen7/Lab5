module Lab5reportQ2Test();
reg [1:0]s;
reg[1:0]I;
wire F;

LabReport5 M1(.s(s),.I(I),.F(F));

initial begin
s[0] = 1'b0;
s[1]= 1'b0;
I[0] = 1'b1;
I[1] = 1'b0;
#100
s[0] = 1'b0;
s[1]= 1'b0;
I[0] = 1'b0;
I[1] = 1'b0;
#100
s[0] = 1'b0;
s[1]= 1'b0;
I[0] = 1'b0;
I[1] = 1'b1;
#100
s[0] = 1'b0;
s[1]= 1'b0;
I[0] = 1'b1;
I[1] = 1'b1;
#100
s[0] = 1'b0;
s[1]= 1'b1;
I[0] = 1'b1;
I[1] = 1'b0;
#100
s[0] = 1'b0;
s[1]= 1'b1;
I[0] = 1'b0;
I[1] = 1'b1;
#100
s[0] = 1'b0;
s[1]= 1'b1;
I[0] = 1'b1;
I[1] = 1'b1;
#100
s[0] = 1'b0;
s[1]= 1'b1;
I[0] = 1'b0;
I[1] = 1'b0;
#100
s[0] = 1'b1;
s[1]= 1'b0;
I[0] = 1'b1;
I[1] = 1'b0;
#100
s[0] = 1'b1;
s[1]= 1'b0;
I[0] = 1'b0;
I[1] = 1'b1;
#100
s[0] = 1'b1;
s[1]= 1'b0;
I[0] = 1'b1;
I[1] = 1'b1;
#100
s[0] = 1'b1;
s[1]= 1'b0;
I[0] = 1'b0;
I[1] = 1'b0;
#100
s[0] = 1'b1;
s[1]= 1'b1;
I[0] = 1'b1;
I[1] = 1'b0;
#100
s[0] = 1'b1;
s[1]= 1'b1;
I[0] = 1'b0;
I[1] = 1'b1;
#100
s[0] = 1'b1;
s[1]= 1'b1;
I[0] = 1'b1;
I[1] = 1'b1;
#100
s[0] = 1'b1;
s[1]= 1'b1;
I[0] = 1'b0;
I[1] = 1'b0;
end
endmodule